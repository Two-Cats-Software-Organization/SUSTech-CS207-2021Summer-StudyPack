`timescale 1ns / 1ps
module project_top_sim(
    );
endmodule
